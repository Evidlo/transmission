.SUBCKT sallenkey n0 out

*define our components
R1  n0 n1 240
R2  n1 in+ 240
RA  in- n4 1K
RB  in- out 10
C1  in+ 0 22pF
C2  n1 out 22pF
X1  in+ in- out n3 0 AD8045

*create vin and power for opamp
VCC n3 0 DC 5.0
VCCvirt n4 0 DC 2.5


.ENDS
